// Course: CSE 401- Computer Architecture
// Term: Winter 2020
// Name: Erika Gutierrez
// ID: 005318270

`timescale 1ns / 1ps

module mem(
   output reg [31:0] data,
   input wire [31:0] addr
   );

   reg [31:0] MEM[0:127];
   integer i;

   initial begin
   MEM[0] <= 'b10001100000000010000000000000001;
   MEM[1] <= 'b10001100000000010000000000000010;
   MEM[2] <= 'b10001100000000010000000000000011;
   MEM[3] <= 'b10000000000000000000000000000000;
   MEM[4] <= 'b10000000000000000000000000000000;
   MEM[5] <= 'b00000000001000100000100000100000;
   MEM[6] <= 'b10000000000000000000000000000000;
   MEM[7] <= 'b10000000000000000000000000000000;
   MEM[8] <= 'b10000000000000000000000000000000;
   MEM[9] <= 'b00000000001000110000100000100000;
   MEM[10] <= 'b10000000000000000000000000000000;
   MEM[11] <= 'b10000000000000000000000000000000;
   MEM[12] <= 'b10000000000000000000000000000000;
   MEM[13] <= 'b00000000001000010000100000100000;
   MEM[14] <= 'b10000000000000000000000000000000;
   MEM[15] <= 'b10000000000000000000000000000000;
   MEM[16] <= 'b10000000000000000000000000000000;
   MEM[17] <= 'b10000000000000000000000000000000;
   MEM[18] <= 'b00000000001000000000100000100000;
   MEM[19] <= 'b10000000000000000000000000000000;
   MEM[20] <= 'b10000000000000000000000000000000;
   MEM[21] <= 'b10000000000000000000000000000000;
   MEM[22] <= 'b10000000000000000000000000000000;
   MEM[23] <= 'b10000000000000000000000000000000;

   // new instructions
   //  MEM[1] <= 'b10001100000000010000000000000000;
   //  MEM[2] <= 'b10001100000001000000000000000001;
   //  MEM[3] <= 'b10000000000000000000000000000000;
   //  MEM[4] <= 'b00000000000000000001000000100000;
   //  MEM[5] <= 'b00000000001000000001100000100000;
   //  MEM[6] <= 'b00010000100000010000000000001110;
   //  MEM[7] <= 'b10000000000000000000000000000000;
   //  MEM[8] <= 'b10000000000000000000000000000000;
   //  MEM[9] <= 'b10000000000000000000000000000000;
   // MEM[10] <= 'b00010000100000000000000000001111;
   // MEM[11] <= 'b10000000000000000000000000000000;
   // MEM[12] <= 'b10000000000000000000000000000000;
   // MEM[13] <= 'b10000000000000000000000000000000;
   // MEM[14] <= 'b00000000010000110001100000100000;
   // MEM[15] <= 'b00000000011000000001000000100000;
   // MEM[16] <= 'b00000000100000010010000000100010;
   // MEM[17] <= 'b00010000000000001111111111110100;
   // MEM[18] <= 'b10000000000000000000000000000000;
   // MEM[19] <= 'b10000000000000000000000000000000;
   // MEM[20] <= 'b10000000000000000000000000000000;
   // MEM[21] <= 'b00000000011000000010100000100000;
   // MEM[22] <= 'b00010000000000000000000000001000;
   // MEM[23] <= 'b10000000000000000000000000000000;
   // MEM[24] <= 'b10000000000000000000000000000000;
   // MEM[25] <= 'b10000000000000000000000000000000;
   // MEM[26] <= 'b00000000010000000010100000100000;
   // MEM[27] <= 'b00010000000000000000000000000011;
   // MEM[28] <= 'b10000000000000000000000000000000;
   // MEM[29] <= 'b10000000000000000000000000000000;
   // MEM[30] <= 'b10000000000000000000000000000000;
   // MEM[31] <= 'b10101100000001010000000000000010;
   // MEM[32] <= 'b10000000000000000000000000000000;
   // MEM[33] <= 'b10000000000000000000000000000000;
   // MEM[34] <= 'b10000000000000000000000000000000;
   // MEM[35] <= 'b10000000000000000000000000000000;
   // MEM[36] <= 'b10000000000000000000000000000000;
   end

   always @(addr) begin
		data <= MEM[addr];
   end
endmodule   //mem
